                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                XXXXXXXX                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        